`include "uvm_macros.svh"

import uvm_pkg::*;

module tb_top;

    initial $display("##--------------TEST STARTED-------------_##");
    final $display("##--------------TEST ENDED--------------##");

    localparam int DATA_WIDTH = 32;
    localparam int SEQ_LENGTH = 32;
    localparam int SHIFT_LEFT = 1;

    logic clk;
    logic arst_n;
    logic serial_in;
    logic we;
    logic [DATA_WIDTH-1:0] parallel_out;   

    ctrl_if ctrl_if();
    data_intf #(DATA_WIDTH) data_if(.clk(clk), .arst_n(arst_n));

    sipo_reg #(
        .DATA_WIDTH(DATA_WIDTH),
        .SHIFT_LEFT(SHIFT_LEFT)
    ) dut (
        .clk(clk),
        .arst_n(arst_n),
        .serial_in(serial_in),
        .we(we),
        .parallel_out(parallel_out)
    );

    assign clk = ctrl_if.clk;
    assign arst_n = ctrl_if.arst_n;
    assign serial_in = data_if.serial_in;
    assign we = data_if.we;
    assign parallel_out = data_if.parallel_out;

    initial begin

        string test;

        if (!$value$plusargs("TEST=%s", test)) begin
            $fatal(1, "No test name provided. Use +TEST=<test_name> to specify a test.");
        end

        $dumpfile("tb_top.vcd");
        $dumpvars(0, tb_top);

        uvm_config_db#(virtual data_intf #(DATA_WIDTH))::set(
            uvm_root::get(), "top", "vif", data_if);
        
        uvm_config_db#(int unsigned)::set(
            uvm_root::get(), "top", "seq_length", SEQ_LENGTH);
        
        uvm_config_db#(int unsigned)::set(
            uvm_root::get(), "top", "shift_left", SHIFT_LEFT);
        

        run_test(test);

        #100 $finish;
    end

endmodule : tb_top